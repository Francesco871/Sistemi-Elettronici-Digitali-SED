library IEEE;
	use IEEE.STD_LOGIC_1164.ALL;

entity HalfAdder is
	Port(
		
	);
end HalfAdder;

architecture Behavioral of HalfAdder is

begin



end Behavioral;
